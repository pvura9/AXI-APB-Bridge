library verilog;
use verilog.vl_types.all;
entity bridgeTop is
end bridgeTop;
