library verilog;
use verilog.vl_types.all;
entity bridgeTop_sv_unit is
end bridgeTop_sv_unit;
